module upper_layer #(
    parameter 
) (
    ports
);
    
endmodule