module process_unit #(
    parameter DATA_WIDTH=8
) ( input clk , rst_n ,
    input  [DATA_WIDTH-1:0] op1,op2,
    output [DATA_WIDTH-1:0] result 
);
    
endmodule